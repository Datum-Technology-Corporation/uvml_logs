// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_LOGS_TDEFS_SV__
`define __UVML_LOGS_TDEFS_SV__


/**
 * 
 */
typedef enum {
   UVML_LOGS_FORMAT_TEXT, ///< 
   UVML_LOGS_FORMAT_JSON, ///< 
   UVML_LOGS_FORMAT_XML , ///< 
   UVML_LOGS_FORMAT_YAML, ///< 
   UVML_LOGS_FORMAT_RAW   ///< 
} uvml_logs_format_enum;


`endif // __UVML_LOGS_TDEFS_SV__
