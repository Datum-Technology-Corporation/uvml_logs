// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVML_LOGS_MACROS_SV__
`define __UVML_LOGS_MACROS_SV__


`define UVML_LOGS_RED   "\033[31m\033[1m"
`define UVML_LOGS_GREEN "\033[32m\033[1m"
`define UVML_LOGS_RESET "\033[0m"


`endif // __UVML_LOGS_MACROS_SV__
