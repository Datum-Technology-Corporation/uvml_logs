// Copyright 2021 Datum Technology Corporation
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


`ifndef __UVME_LOGS_ST_CONSTANTS_SV__
`define __UVME_LOGS_ST_CONSTANTS_SV__





`endif // __UVME_LOGS_ST_CONSTANTS_SV__
